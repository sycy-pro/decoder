module brute_force(
    input clk,
    input rst,
    input ena,
    input start,
    input [63:0] data,
    
    output [47:0] key_out,
    output valid,
    output rdy
);

localparam DICT4_SIZE = 2500;

localparam bit [31:0] DICT4 [DICT4_SIZE-1:0]= '{
32'h77656573,
32'h77656570,
32'h7765656e,
32'h7765656c,
32'h77656473,
32'h77656273,
32'h7765616e,
32'h7765616c,
32'h77617879,
32'h77617679,
32'h77617474,
32'h77617374,
32'h77617370,
32'h77617274,
32'h77617270,
32'h77617265,
32'h77616e73,
32'h77616e65,
32'h77616e64,
32'h77616c69,
32'h77616c65,
32'h7761696c,
32'h77616966,
32'h77616773,
32'h77616674,
32'h77616473,
32'h77616469,
32'h77616465,
32'h7761636b,
32'h766f7773,
32'h766f6c65,
32'h76697661,
32'h76697461,
32'h76697365,
32'h76696f6c,
32'h76696e6f,
32'h76696d73,
32'h76696c6c,
32'h76696c65,
32'h76696573,
32'h76696564,
32'h76696473,
32'h7669616c,
32'h76657473,
32'h7665746f,
32'h76657274,
32'h76656e64,
32'h76656e61,
32'h76656c64,
32'h7665696c,
32'h76656573,
32'h76656572,
32'h76656570,
32'h7665616c,
32'h76617473,
32'h76617365,
32'h76617361,
32'h76616e73,
32'h76616e65,
32'h76616d70,
32'h76616c65,
32'h7661696e,
32'h7661696c,
32'h76616373,
32'h75726e73,
32'h75726963,
32'h75726561,
32'h7570646f,
32'h756e646f,
32'h756d7073,
32'h756d6d61,
32'h756c6e61,
32'h75646f6e,
32'h7479726f,
32'h7479706f,
32'h74796b65,
32'h74776f73,
32'h74776974,
32'h74776967,
32'h74776565,
32'h74757475,
32'h74757473,
32'h7475736b,
32'h74757368,
32'h7475726b,
32'h74757264,
32'h74756d73,
32'h74756c65,
32'h74756773,
32'h74756674,
32'h74756666,
32'h74756661,
32'h7475636b,
32'h74756273,
32'h74756261,
32'h74736172,
32'h74727565,
32'h74726f74,
32'h74726f64,
32'h74726967,
32'h74726579,
32'h7472656b,
32'h7472616d,
32'h746f7773,
32'h746f7574,
32'h746f7473,
32'h746f7465,
32'h746f7279,
32'h746f7274,
32'h746f7272,
32'h746f7265,
32'h746f7263,
32'h746f706f,
32'h746f7069,
32'h746f6f74,
32'h746f6f6e,
32'h746f6e79,
32'h746f6e67,
32'h746f6d65,
32'h746f6c65,
32'h746f6b65,
32'h746f696c,
32'h746f6761,
32'h746f6675,
32'h746f6666,
32'h746f6564,
32'h746f6279,
32'h746f6164,
32'h74697069,
32'h74696e74,
32'h74696e73,
32'h74696e67,
32'h74696e65,
32'h74696c74,
32'h74696b69,
32'h74696666,
32'h74696479,
32'h74696373,
32'h7469616e,
32'h74687567,
32'h74687564,
32'h7468726f,
32'h74686577,
32'h74686177,
32'h7465726e,
32'h74656c65,
32'h74656666,
32'h74656573,
32'h7465656d,
32'h74656174,
32'h74656173,
32'h7465616c,
32'h7465616b,
32'h74617861,
32'h74617574,
32'h74617274,
32'h74617273,
32'h74617270,
32'h7461726f,
32'h7461726e,
32'h74617265,
32'h74617073,
32'h74617061,
32'h74616e73,
32'h74616e67,
32'h74616d70,
32'h74616d65,
32'h74616c63,
32'h74616374,
32'h7461636f,
32'h7461636b,
32'h74616368,
32'h74616275,
32'h7377756d,
32'h73776967,
32'h73776179,
32'h73776174,
32'h7377616e,
32'h7377616d,
32'h73776167,
32'h73776162,
32'h73757373,
32'h73757261,
32'h73757073,
32'h73756e73,
32'h73756e6b,
32'h73756e67,
32'h73756d73,
32'h73756d70,
32'h73756d6f,
32'h73756c6b,
32'h73756574,
32'h73756573,
32'h73756273,
32'h73747965,
32'h7374756e,
32'h73747564,
32'h73747562,
32'h73746f77,
32'h73746577,
32'h73746167,
32'h73746162,
32'h73707572,
32'h7370756e,
32'h73707564,
32'h73707279,
32'h73706974,
32'h73706963,
32'h73706577,
32'h73706564,
32'h7370617a,
32'h73706179,
32'h73706174,
32'h73706173,
32'h73706172,
32'h736f7961,
32'h736f7773,
32'h736f776e,
32'h736f756b,
32'h736f7473,
32'h736f7261,
32'h736f7073,
32'h736f6f74,
32'h736f6d61,
32'h736f6473,
32'h736f636b,
32'h736f6361,
32'h736f6273,
32'h736f6261,
32'h736f6172,
32'h736e7567,
32'h736e7562,
32'h736e6f74,
32'h736e6f67,
32'h736e6f62,
32'h736e6974,
32'h736e6970,
32'h736e6167,
32'h736d7574,
32'h736d7567,
32'h736d6f67,
32'h736c7572,
32'h736c756d,
32'h736c7567,
32'h736c6f70,
32'h736c6f67,
32'h736c6f65,
32'h736c6f62,
32'h736c6974,
32'h736c6964,
32'h736c6577,
32'h736c6564,
32'h736c6179,
32'h736c6177,
32'h736c6174,
32'h736c6170,
32'h736c616d,
32'h736c6167,
32'h736c6162,
32'h736b7561,
32'h736b6974,
32'h736b6973,
32'h736b696d,
32'h736b6964,
32'h736b6577,
32'h736b6567,
32'h73697273,
32'h73697265,
32'h73697073,
32'h73696e65,
32'h73696c74,
32'h73696c6f,
32'h73696c6c,
32'h73696b61,
32'h73696768,
32'h73696674,
32'h73696273,
32'h7368756e,
32'h7368756c,
32'h73686f6f,
32'h73686f64,
32'h73686976,
32'h7368696e,
32'h7368696d,
32'h73686577,
32'h7368616d,
32'h73686168,
32'h73686167,
32'h73686164,
32'h73657773,
32'h7365776e,
32'h73657474,
32'h73657461,
32'h73657266,
32'h73657265,
32'h73657074,
32'h73656d69,
32'h73656572,
32'h73656570,
32'h73656374,
32'h73656172,
32'h7363756d,
32'h73637564,
32'h73636f77,
32'h73636f74,
32'h73636174,
32'h73636172,
32'h73636164,
32'h73636162,
32'h73617773,
32'h7361776e,
32'h73617469,
32'h73617465,
32'h73617373,
32'h73617368,
32'h73617269,
32'h73617073,
32'h73616e6b,
32'h73616e65,
32'h73616b69,
32'h73616773,
32'h7361676f,
32'h73616373,
32'h7361636b,
32'h72757473,
32'h72757468,
32'h72757365,
32'h72756e74,
32'h72756e67,
32'h72756e65,
32'h72756d73,
32'h72756d70,
32'h72756773,
32'h72756666,
32'h72756573,
32'h72756564,
32'h7275636b,
32'h72756279,
32'h72756273,
32'h72756265,
32'h726f7665,
32'h726f7578,
32'h726f7574,
32'h726f7473,
32'h726f746f,
32'h726f7469,
32'h726f7465,
32'h726f7461,
32'h726f7379,
32'h726f7079,
32'h726f6f73,
32'h726f6f6b,
32'h726f6f64,
32'h726f6d73,
32'h726f6d70,
32'h726f696c,
32'h726f6573,
32'h726f6273,
32'h726f6265,
32'h726f6172,
32'h726f616e,
32'h726f616d,
32'h7269747a,
32'h72697465,
32'h72697073,
32'h72696f74,
32'h72696e6b,
32'h72696e64,
32'h72696d73,
32'h72696d65,
32'h72696c6c,
32'h72696c65,
32'h72696773,
32'h72696674,
32'h72696666,
32'h72696665,
32'h72696473,
32'h72686561,
32'h72657465,
32'h72657070,
32'h7265706f,
32'h72656e64,
32'h72656d73,
32'h7265696e,
32'h72656673,
32'h7265656b,
32'h72656564,
32'h7265646f,
32'h7265616d,
32'h72617a7a,
32'h72617a65,
32'h72617665,
32'h72617468,
32'h72617370,
32'h72617074,
32'h72617073,
32'h72616e74,
32'h72616e67,
32'h72616d73,
32'h72616d69,
32'h72616c65,
32'h72616b75,
32'h72616b69,
32'h72616b65,
32'h72616a61,
32'h72616773,
32'h72616761,
32'h72616674,
32'h72616473,
32'h72616379,
32'h71756970,
32'h71756964,
32'h71756179,
32'h7079726f,
32'h70797265,
32'h7075747a,
32'h70757474,
32'h70757373,
32'h70757272,
32'h7075726c,
32'h70757269,
32'h70757073,
32'h70757061,
32'h70756e79,
32'h70756e74,
32'h70756e73,
32'h70756d61,
32'h70756c70,
32'h70756b65,
32'h70756a61,
32'h70756773,
32'h70756666,
32'h70756473,
32'h70736973,
32'h70726f77,
32'h70726f6d,
32'h70726f67,
32'h70726f66,
32'h70726f64,
32'h70726f62,
32'h7072696d,
32'h70726967,
32'h7072657a,
32'h7072616d,
32'h706f7879,
32'h706f7574,
32'h706f7566,
32'h706f7379,
32'h706f7368,
32'h706f7265,
32'h706f6f70,
32'h706f6f66,
32'h706f6e79,
32'h706f6e67,
32'h706f6e65,
32'h706f6d70,
32'h706f6d65,
32'h706f6c79,
32'h706f6c73,
32'h706f6b79,
32'h706f6b65,
32'h706f6473,
32'h706f636b,
32'h706c756d,
32'h706c6f79,
32'h706c6f77,
32'h706c6f70,
32'h706c6f64,
32'h706c6578,
32'h706c6564,
32'h706c6562,
32'h706c6174,
32'h70697879,
32'h70697479,
32'h70697473,
32'h70697468,
32'h70697461,
32'h70697373,
32'h70697368,
32'h70697061,
32'h70696f6e,
32'h70696e74,
32'h70696e67,
32'h70696d70,
32'h70696b65,
32'h70696b61,
32'h70696573,
32'h70696564,
32'h70696365,
32'h70696361,
32'h70686973,
32'h70686577,
32'h70657773,
32'h7065736f,
32'h70657276,
32'h70657274,
32'h70657270,
32'h7065726d,
32'h7065726b,
32'h70657269,
32'h7065706f,
32'h70656f6e,
32'h70656e74,
32'h70656c74,
32'h70656773,
32'h70656573,
32'h70656570,
32'h7065656b,
32'h70656564,
32'h70656473,
32'h70656373,
32'h7065636b,
32'h70656174,
32'h70656172,
32'h7065616c,
32'h70617773,
32'h7061776e,
32'h70617665,
32'h70617473,
32'h70617465,
32'h70617273,
32'h70617265,
32'h70617261,
32'h70617073,
32'h70617061,
32'h70616e74,
32'h70616e67,
32'h70616c73,
32'h70616c70,
32'h70616c6c,
32'h7061696c,
32'h70616374,
32'h6f776c73,
32'h6f776573,
32'h6f76756d,
32'h6f76616c,
32'h6f757a6f,
32'h6f757374,
32'h6f756368,
32'h6f74746f,
32'h6f746963,
32'h6f727a6f,
32'h6f727978,
32'h6f726779,
32'h6f726573,
32'h6f72646f,
32'h6f726361,
32'h6f726273,
32'h6f707573,
32'h6f707473,
32'h6f70616c,
32'h6f6f7a79,
32'h6f6f7a65,
32'h6f6f7073,
32'h6f6e7978,
32'h6f6e7573,
32'h6f6d6974,
32'h6f6d656e,
32'h6f6c6c61,
32'h6f6c656f,
32'h6f6c6479,
32'h6f6c6473,
32'h6f6b7261,
32'h6f696e6b,
32'h6f677265,
32'h6f676c65,
32'h6f676565,
32'h6f646573,
32'h6f626f65,
32'h6f626974,
32'h6f617273,
32'h6f616b79,
32'h6f616b73,
32'h6f616673,
32'h6e756e73,
32'h6e756d62,
32'h6e756b65,
32'h6e756273,
32'h6e6f7661,
32'h6e6f7573,
32'h6e6f756e,
32'h6e6f7379,
32'h6e6f7368,
32'h6e6f7269,
32'h6e6f6f6b,
32'h6e6f6d65,
32'h6e6f6972,
32'h6e6f656c,
32'h6e6f6473,
32'h6e6f636b,
32'h6e6f6273,
32'h6e697465,
32'h6e697073,
32'h6e696768,
32'h6e69636b,
32'h6e696273,
32'h6e657774,
32'h6e657373,
32'h6e657264,
32'h6e656f6e,
32'h6e656e65,
32'h6e65656d,
32'h6e656170,
32'h6e617973,
32'h6e617665,
32'h6e617279,
32'h6e617264,
32'h6e617263,
32'h6e617073,
32'h6e617065,
32'h6e617061,
32'h6e616e73,
32'h6e616e61,
32'h6e616773,
32'h6e616666,
32'h6e616273,
32'h6e616265,
32'h6e61616e,
32'h6d757474,
32'h6d757465,
32'h6d757373,
32'h6d75736b,
32'h6d757368,
32'h6d757365,
32'h6d75726b,
32'h6d756f6e,
32'h6d756e67,
32'h6d756d73,
32'h6d756c6c,
32'h6d756c65,
32'h6d756773,
32'h6d756666,
32'h6d756473,
32'h6d75636b,
32'h6d6f7773,
32'h6d6f7468,
32'h6d6f7465,
32'h6d6f7373,
32'h6d6f7368,
32'h6d6f726e,
32'h6d6f7073,
32'h6d6f7065,
32'h6d6f6f74,
32'h6d6f6f73,
32'h6d6f6f72,
32'h6d6f6f6b,
32'h6d6f6e6f,
32'h6d6f6e6b,
32'h6d6f6c74,
32'h6d6f6c6c,
32'h6d6f6c65,
32'h6d6f6c61,
32'h6d6f6a6f,
32'h6d6f636b,
32'h6d6f6273,
32'h6d6f6174,
32'h6d6f616e,
32'h6d697474,
32'h6d697465,
32'h6d69736f,
32'h6d697365,
32'h6d697279,
32'h6d697265,
32'h6d696e78,
32'h6d696e6b,
32'h6d696e61,
32'h6d696d65,
32'h6d696b65,
32'h6d69656e,
32'h6d696473,
32'h6d696373,
32'h6d696361,
32'h6d657a65,
32'h6d657773,
32'h6d65776c,
32'h6d657465,
32'h6d657461,
32'h6d657361,
32'h6d656f77,
32'h6d656e64,
32'h6d656d6f,
32'h6d656c64,
32'h6d65656b,
32'h6d656164,
32'h6d617a79,
32'h6d617a65,
32'h6d61796f,
32'h6d617961,
32'h6d617869,
32'h6d617773,
32'h6d61756c,
32'h6d617374,
32'h6d617368,
32'h6d617361,
32'h6d617274,
32'h6d617273,
32'h6d61726c,
32'h6d617265,
32'h6d616e65,
32'h6d616c74,
32'h6d616b6f,
32'h6d616b69,
32'h6d61696d,
32'h6d616964,
32'h6d616773,
32'h6d616769,
32'h6d616765,
32'h6d616373,
32'h6d61636b,
32'h6d616368,
32'h6d616365,
32'h6c797365,
32'h6c797265,
32'h6c796e78,
32'h6c757673,
32'h6c757465,
32'h6c757374,
32'h6c75726b,
32'h6c757265,
32'h6c756e65,
32'h6c756c6c,
32'h6c756773,
32'h6c756765,
32'h6c756666,
32'h6c756265,
32'h6c756175,
32'h6c6f7773,
32'h6c6f7574,
32'h6c6f7468,
32'h6c6f7265,
32'h6c6f7073,
32'h6c6f7065,
32'h6c6f6f74,
32'h6c6f6f73,
32'h6c6f6f6e,
32'h6c6f6f6d,
32'h6c6f6c6c,
32'h6c6f696e,
32'h6c6f6765,
32'h6c6f6465,
32'h6c6f636f,
32'h6c6f6368,
32'h6c6f6273,
32'h6c6f6265,
32'h6c6f616d,
32'h6c6f6166,
32'h6c697465,
32'h6c697370,
32'h6c697261,
32'h6c696e74,
32'h6c696e67,
32'h6c696d70,
32'h6c696d6f,
32'h6c696d6e,
32'h6c696d61,
32'h6c696c79,
32'h6c696c74,
32'h6c696575,
32'h6c696572,
32'h6c69656e,
32'h6c696564,
32'h6c696473,
32'h6c69636b,
32'h6c696365,
32'h6c696273,
32'h6c696172,
32'h6c657973,
32'h6c657764,
32'h6c657679,
32'h6c657374,
32'h6c656e74,
32'h6c656973,
32'h6c656574,
32'h6c656572,
32'h6c65656b,
32'h6c656173,
32'h6c617a65,
32'h6c617665,
32'h6c617564,
32'h6c617473,
32'h6c617468,
32'h6c617373,
32'h6c617368,
32'h6c61726b,
32'h6c617264,
32'h6c617073,
32'h6c616d73,
32'h6c616d65,
32'h6c616d61,
32'h6c616b68,
32'h6c616972,
32'h6c61696e,
32'h6c616773,
32'h6c616473,
32'h6c616379,
32'h6b756475,
32'h6b6f746f,
32'h6b6f7261,
32'h6b6f6f6b,
32'h6b6f6c61,
32'h6b6f6a69,
32'h6b6f686c,
32'h6b6f616e,
32'h6b697769,
32'h6b697661,
32'h6b697468,
32'h6b697465,
32'h6b697073,
32'h6b696c74,
32'h6b696c6f,
32'h6b696c6e,
32'h6b686174,
32'h6b68616e,
32'h6b65746f,
32'h6b657266,
32'h6b657262,
32'h6b656c70,
32'h6b656773,
32'h6b65656c,
32'h6b617661,
32'h6b617461,
32'h6b617274,
32'h6b616d69,
32'h6b616c65,
32'h6b616b61,
32'h6a757473,
32'h6a757465,
32'h6a756b65,
32'h6a756a75,
32'h6a756773,
32'h6a756479,
32'h6a75646f,
32'h6a6f7973,
32'h6a6f776c,
32'h6a6f7473,
32'h6a6f7368,
32'h6a6f6c74,
32'h6a6f686e,
32'h6a6f6773,
32'h6a6f6579,
32'h6a6f636b,
32'h6a697665,
32'h6a696e78,
32'h6a696e6e,
32'h6a696e6b,
32'h6a696c74,
32'h6a696773,
32'h6a696273,
32'h6a696265,
32'h6a657374,
32'h6a65726b,
32'h6a656c6c,
32'h6a656665,
32'h6a65657a,
32'h6a656572,
32'h6a65616e,
32'h6a617973,
32'h6a617773,
32'h6a617661,
32'h6a617065,
32'h6a616d73,
32'h6a616d62,
32'h6a616b65,
32'h6a616465,
32'h6a616273,
32'h69746368,
32'h69736d73,
32'h69726b73,
32'h69726973,
32'h696f7461,
32'h696e6e73,
32'h696e6b79,
32'h696e6b73,
32'h696d7073,
32'h696d616d,
32'h696c6c73,
32'h696b6f6e,
32'h696b6174,
32'h69666679,
32'h69646f6c,
32'h69646c79,
32'h69636b79,
32'h69636573,
32'h69636564,
32'h69626973,
32'h69626578,
32'h6879706f,
32'h68796d6e,
32'h68757473,
32'h6875736b,
32'h68757368,
32'h6875726c,
32'h68756e6b,
32'h68756d73,
32'h68756d70,
32'h68756c6b,
32'h68756c61,
32'h68756773,
32'h68756666,
32'h68756573,
32'h68756564,
32'h6875636b,
32'h686f776c,
32'h686f7665,
32'h686f7261,
32'h686f7073,
32'h686f6f74,
32'h686f6f70,
32'h686f6f66,
32'h686f6e6b,
32'h686f6e67,
32'h686f6e65,
32'h686f6c74,
32'h686f6c6f,
32'h686f6773,
32'h686f6573,
32'h686f6564,
32'h686f636b,
32'h686f626f,
32'h686f6178,
32'h686f6172,
32'h68697961,
32'h68697665,
32'h68697373,
32'h68696e64,
32'h68696c74,
32'h68696564,
32'h6869636b,
32'h68657773,
32'h6865776e,
32'h68656e73,
32'h68656d73,
32'h68656d65,
32'h68656c6f,
32'h68656c6d,
32'h68656972,
32'h68656674,
32'h68656564,
32'h68656170,
32'h68617a79,
32'h68617a65,
32'h68617973,
32'h68617773,
32'h6861776b,
32'h6861756c,
32'h68617370,
32'h68617274,
32'h68617270,
32'h6861726b,
32'h68617265,
32'h68617073,
32'h68616e6b,
32'h68616d73,
32'h68616c74,
32'h68616b65,
32'h68616a6a,
32'h6861696c,
32'h68616773,
32'h68616674,
32'h6779726f,
32'h67797265,
32'h67796d73,
32'h67757473,
32'h67757374,
32'h67757368,
32'h67756e6b,
32'h67756d73,
32'h67756c70,
32'h67756c6c,
32'h67756666,
32'h67756172,
32'h67727565,
32'h67727562,
32'h67726f67,
32'h67726974,
32'h6772696e,
32'h6772696d,
32'h67726565,
32'h6772616e,
32'h6772616d,
32'h67726164,
32'h676f7973,
32'h676f7574,
32'h676f7468,
32'h676f7368,
32'h676f7279,
32'h676f7265,
32'h676f6f73,
32'h676f6f70,
32'h676f6f6e,
32'h676f6f6b,
32'h676f6f66,
32'h676f6e67,
32'h676f6572,
32'h676f6279,
32'h676f6273,
32'h676f6164,
32'h676e7573,
32'h676e6177,
32'h676e6174,
32'h676e6172,
32'h676c7574,
32'h676c756d,
32'h676c7567,
32'h676c6f70,
32'h676c6f6d,
32'h676c6f62,
32'h676c6962,
32'h676c6961,
32'h676c656e,
32'h676c6565,
32'h676c616d,
32'h67697473,
32'h67697465,
32'h67697374,
32'h67697274,
32'h67697264,
32'h67696e73,
32'h67696d70,
32'h67696c74,
32'h67696c6c,
32'h67696c64,
32'h67696773,
32'h67696265,
32'h67686565,
32'h67686174,
32'h67657461,
32'h6765726d,
32'h67656e75,
32'h67656e74,
32'h67656e73,
32'h67656c74,
32'h67656c73,
32'h67656573,
32'h6765656b,
32'h67617973,
32'h67617770,
32'h6761776b,
32'h67617370,
32'h67617368,
32'h67617262,
32'h67617065,
32'h67616f6c,
32'h67616d73,
32'h67616c73,
32'h67616c6c,
32'h67616c65,
32'h67616c61,
32'h67616974,
32'h67616773,
32'h67616765,
32'h67616666,
32'h66757a7a,
32'h6675747a,
32'h66757373,
32'h66757273,
32'h6675726c,
32'h66756e6b,
32'h66756d65,
32'h66756775,
32'h66726967,
32'h66726574,
32'h66726179,
32'h66726174,
32'h66726167,
32'h666f7879,
32'h666f776c,
32'h666f756c,
32'h666f7265,
32'h666f7264,
32'h666f7073,
32'h666f6779,
32'h666f6773,
32'h666f6573,
32'h666f6369,
32'h666f6273,
32'h666f616c,
32'h666c7578,
32'h666c7573,
32'h666c7565,
32'h666c7562,
32'h666c6f70,
32'h666c6f67,
32'h666c6f65,
32'h666c6f63,
32'h666c6974,
32'h666c6565,
32'h666c6561,
32'h666c6179,
32'h666c6178,
32'h666c6177,
32'h666c6170,
32'h666c616e,
32'h666c616d,
32'h666c616b,
32'h666c6162,
32'h66697a7a,
32'h66697273,
32'h66696e73,
32'h66696e6b,
32'h66696c6f,
32'h66696773,
32'h66696665,
32'h66696566,
32'h66696273,
32'h66696174,
32'h66657564,
32'h66657465,
32'h66657461,
32'h66657374,
32'h66657373,
32'h6665726e,
32'h66656e73,
32'h66656e64,
32'h6665636b,
32'h66617a65,
32'h6661776e,
32'h66617665,
32'h66617661,
32'h6661756e,
32'h66617274,
32'h6661726f,
32'h66616e67,
32'h6661696e,
32'h66616473,
32'h6661646f,
32'h66616273,
32'h65796564,
32'h6578706f,
32'h65786f6e,
32'h65786563,
32'h65776573,
32'h65776572,
32'h65766573,
32'h65746368,
32'h65746173,
32'h65727576,
32'h65727273,
32'h65726773,
32'h65726173,
32'h65706565,
32'h656f6e73,
32'h656e7679,
32'h656d7573,
32'h656d6d79,
32'h656d6974,
32'h656d6972,
32'h656d6963,
32'h656c6d73,
32'h656c6c73,
32'h656c6b73,
32'h656c616e,
32'h656b6573,
32'h65676f73,
32'h65676779,
32'h65656c73,
32'h65646779,
32'h65646479,
32'h65637275,
32'h65626273,
32'h65617665,
32'h64796b65,
32'h64796573,
32'h64796572,
32'h64796564,
32'h64796164,
32'h6475736b,
32'h64757261,
32'h64757065,
32'h64756f73,
32'h64756e73,
32'h64756e6b,
32'h64756e67,
32'h64756e65,
32'h64756c79,
32'h64756773,
32'h64756666,
32'h64756574,
32'h64756573,
32'h6475656c,
32'h64756473,
32'h64756273,
32'h64727973,
32'h64726970,
32'h64726179,
32'h6472616d,
32'h64726162,
32'h646f7a79,
32'h646f7a65,
32'h646f7879,
32'h646f7665,
32'h646f7572,
32'h646f7468,
32'h646f7465,
32'h646f7361,
32'h646f7279,
32'h646f726d,
32'h646f726b,
32'h646f7065,
32'h646f6e67,
32'h646f6c74,
32'h646f6c65,
32'h646f6a6f,
32'h646f6765,
32'h646f6666,
32'h646f6572,
32'h646f646f,
32'h64697661,
32'h64697373,
32'h64697265,
32'h64697073,
32'h64696e74,
32'h64696e6f,
32'h64696e6b,
32'h64696e67,
32'h64696e65,
32'h64696d73,
32'h64696d65,
32'h64696c6c,
32'h64696b65,
32'h64696773,
32'h64686f77,
32'h6468616c,
32'h64657779,
32'h64657773,
32'h6465726d,
32'h64656e74,
32'h64656e73,
32'h64656c74,
32'h64656c6c,
32'h64656c69,
32'h64656b65,
32'h64656679,
32'h64656674,
32'h6465656d,
32'h6465616e,
32'h64617a65,
32'h64617562,
32'h64617274,
32'h6461726e,
32'h64616e6b,
32'h64616d73,
32'h64616d65,
32'h64616c65,
32'h64616973,
32'h64616674,
32'h64616473,
32'h6461646f,
32'h64616461,
32'h64616365,
32'h64616273,
32'h637a6172,
32'h63797374,
32'h6379616e,
32'h63757373,
32'h63757370,
32'h63757274,
32'h63757273,
32'h6375726c,
32'h63757264,
32'h63757262,
32'h63756c6d,
32'h63756c6c,
32'h63756666,
32'h63756564,
32'h63756473,
32'h63727578,
32'h63727573,
32'h63727564,
32'h63726f77,
32'h63726f63,
32'h63726974,
32'h63726962,
32'h63726177,
32'h6372616d,
32'h63726167,
32'h636f776c,
32'h636f7570,
32'h636f7473,
32'h636f7465,
32'h636f7379,
32'h636f7368,
32'h636f726d,
32'h636f726b,
32'h636f6f74,
32'h636f6f73,
32'h636f6f70,
32'h636f6e6e,
32'h636f6e6b,
32'h636f6d70,
32'h636f6d62,
32'h636f6d61,
32'h636f6c74,
32'h636f6c65,
32'h636f6c61,
32'h636f6972,
32'h636f6966,
32'h636f686f,
32'h636f6773,
32'h636f6564,
32'h636f6473,
32'h636f6461,
32'h636f636f,
32'h636f6361,
32'h636f6273,
32'h636f6178,
32'h636c6f74,
32'h636c6f70,
32'h636c6f67,
32'h636c6f64,
32'h636c6566,
32'h636c6177,
32'h636c6170,
32'h636c616d,
32'h636c6164,
32'h63697465,
32'h6369616f,
32'h6368756d,
32'h63687567,
32'h63687562,
32'h63686f77,
32'h63686974,
32'h63686172,
32'h63686170,
32'h63686169,
32'h63686164,
32'h63657373,
32'h63656c74,
32'h63656c73,
32'h63656465,
32'h63617973,
32'h63617773,
32'h63617679,
32'h63617661,
32'h6361756c,
32'h6361736b,
32'h63617272,
32'h63617270,
32'h6361706f,
32'h63617065,
32'h63616d73,
32'h63616d6f,
32'h63616d69,
32'h63616666,
32'h63616473,
32'h63616273,
32'h62797465,
32'h62797265,
32'h62796573,
32'h62757a7a,
32'h62757374,
32'h62757373,
32'h6275736b,
32'h62757279,
32'h62757272,
32'h62757270,
32'h6275726c,
32'h62757267,
32'h62757262,
32'h62756f79,
32'h62756e74,
32'h62756e73,
32'h62756e6b,
32'h62756e67,
32'h62756e64,
32'h62756d73,
32'h62756666,
32'h62726f77,
32'h62726f73,
32'h62726974,
32'h62726973,
32'h6272696f,
32'h6272696d,
32'h62726967,
32'h62726965,
32'h62726564,
32'h62726179,
32'h62726174,
32'h62726173,
32'h6272616e,
32'h62726167,
32'h62726164,
32'h626f7a6f,
32'h626f796f,
32'h626f7879,
32'h626f7773,
32'h626f7473,
32'h626f6f73,
32'h626f6f72,
32'h626f6f6e,
32'h626f6f62,
32'h626f6e79,
32'h626f6e6b,
32'h626f6e67,
32'h626f6c6f,
32'h626f6c6c,
32'h626f6c65,
32'h626f6c61,
32'h626f6779,
32'h626f6773,
32'h626f6473,
32'h626f6465,
32'h626f6273,
32'h626f6173,
32'h626f6172,
32'h626c7572,
32'h626c6f74,
32'h626c6f63,
32'h626c6f62,
32'h626c6970,
32'h626c6564,
32'h626c6562,
32'h626c6162,
32'h62696f73,
32'h62696e74,
32'h62696c6b,
32'h62696c65,
32'h62696666,
32'h62696572,
32'h62696465,
32'h62696273,
32'h62696262,
32'h62657973,
32'h62657679,
32'h62657473,
32'h6265726d,
32'h62657267,
32'h62656773,
32'h62656574,
32'h62656570,
32'h6265636b,
32'h62656175,
32'h6265616b,
32'h62617973,
32'h6261776c,
32'h62617564,
32'h62617474,
32'h62617374,
32'h6261736b,
32'h62617368,
32'h62617266,
32'h62617264,
32'h62617262,
32'h62616e73,
32'h62616e65,
32'h62616c6d,
32'h62616c6b,
32'h62616c65,
32'h62616c64,
32'h62616874,
32'h62616473,
32'h62616465,
32'h62616368,
32'h62616265,
32'h62616261,
32'h61786f6e,
32'h6178696c,
32'h61786573,
32'h6178656c,
32'h61786564,
32'h61777279,
32'h61776c73,
32'h61776573,
32'h61776564,
32'h61766f77,
32'h61766572,
32'h61736879,
32'h6172796c,
32'h6172756d,
32'h61727479,
32'h61727365,
32'h61726b73,
32'h6172696c,
32'h61726964,
32'h61726961,
32'h61726373,
32'h61717561,
32'h61707365,
32'h61706578,
32'h61706573,
32'h616e6f6e,
32'h616e6e61,
32'h616e6b68,
32'h616e6577,
32'h616e6473,
32'h616d796c,
32'h616d6f6b,
32'h616d626f,
32'h616c756d,
32'h616c746f,
32'h616c6f65,
32'h616c6d73,
32'h616c6761,
32'h616c6573,
32'h616c6172,
32'h616a6172,
32'h61697279,
32'h61697273,
32'h61696c73,
32'h61696465,
32'h6168656d,
32'h61677565,
32'h61676f67,
32'h61676172,
32'h6166726f,
32'h61666172,
32'h61656f6e,
32'h61647a65,
32'h61646974,
32'h61636d65,
32'h61636879,
32'h61636865,
32'h61636573,
32'h61636564,
32'h61636169,
32'h61627574,
32'h61626c79,
32'h61626574,
32'h61626564,
32'h7a6f6f6d,
32'h7a696e63,
32'h7961726e,
32'h776f726d,
32'h776f6f6c,
32'h776f6c66,
32'h776f6b65,
32'h77697065,
32'h77656564,
32'h77617279,
32'h7761726e,
32'h77617264,
32'h766f6c74,
32'h766f6964,
32'h76696e65,
32'h76696265,
32'h76657374,
32'h76657262,
32'h76656e74,
32'h7665696e,
32'h75726765,
32'h74797265,
32'h74757266,
32'h74756e61,
32'h7472696f,
32'h7472696d,
32'h74726179,
32'h74726170,
32'h746f7373,
32'h746f726e,
32'h746f7073,
32'h746f6d62,
32'h746f6c6c,
32'h746f6573,
32'h74696573,
32'h74696465,
32'h7469636b,
32'h74687275,
32'h74686565,
32'h74656d70,
32'h74656172,
32'h74617869,
32'h74616273,
32'h7377696d,
32'h73776170,
32'h73757266,
32'h73756564,
32'h7375636b,
32'h73746174,
32'h7370696e,
32'h73706563,
32'h7370616e,
32'h736f7572,
32'h736f7265,
32'h736f6661,
32'h736f616b,
32'h736e6170,
32'h736c6970,
32'h736c696d,
32'h73696e73,
32'h73696e6b,
32'h73696c6b,
32'h73686564,
32'h73657879,
32'h73656173,
32'h7365616d,
32'h7363616d,
32'h73616e67,
32'h7361696c,
32'h73616765,
32'h73616761,
32'h72757374,
32'h72757368,
32'h7275696e,
32'h72756465,
32'h726f6473,
32'h726f6465,
32'h72697065,
32'h72696273,
32'h72657073,
32'h7265656c,
32'h72656566,
32'h72656170,
32'h72617973,
32'h72617473,
32'h72617368,
32'h72617065,
32'h72616d70,
32'h72616964,
32'h72616765,
32'h7175697a,
32'h71756164,
32'h70756e6b,
32'h7075636b,
32'h70756273,
32'h70726f70,
32'h70726579,
32'h706f7473,
32'h706f7365,
32'h706f726e,
32'h706f726b,
32'h706f7073,
32'h706f7065,
32'h706f6e64,
32'h706f6c6f,
32'h706f6574,
32'h706f656d,
32'h706c6561,
32'h70696e65,
32'h70696c6c,
32'h70696c65,
32'h70696773,
32'h70696572,
32'h70696373,
32'h70657374,
32'h70656e73,
32'h70656572,
32'h7065656c,
32'h70656173,
32'h70616e73,
32'h70616e65,
32'h70616c65,
32'h6f776564,
32'h6f757473,
32'h6f757273,
32'h6f696c79,
32'h6f646f72,
32'h6f626579,
32'h6f617473,
32'h6f617468,
32'h6e756c6c,
32'h6e756465,
32'h6e6f726d,
32'h6e6f7065,
32'h6e6f6f6e,
32'h6e657473,
32'h6e657374,
32'h6d797468,
32'h6d6f6d73,
32'h6d6f6c64,
32'h6d6f6473,
32'h6d697374,
32'h6d696e74,
32'h6d696365,
32'h6d656c74,
32'h6d656761,
32'h6d617473,
32'h6d617465,
32'h6d616e73,
32'h6d616d61,
32'h6c757368,
32'h6c756e67,
32'h6c756d70,
32'h6c6f7564,
32'h6c6f6e65,
32'h6c6f6773,
32'h6c6f6674,
32'h6c696f6e,
32'h6c696d65,
32'h6c696d62,
32'h6c656e64,
32'h6c656170,
32'h6c65616e,
32'h6c65616b,
32'h6c617a79,
32'h6c617973,
32'h6c617661,
32'h6c616d70,
32'h6c616d62,
32'h6c616365,
32'h6c616273,
32'h6b6e6f74,
32'h6b6e6f62,
32'h6b6e6974,
32'h6b697373,
32'h6a756e6b,
32'h6a657473,
32'h6a656570,
32'h6a617273,
32'h6a61636b,
32'h69736c65,
32'h696f6e73,
32'h69646c65,
32'h68797065,
32'h68756e74,
32'h68756e67,
32'h68756c6c,
32'h68756273,
32'h686f726e,
32'h686f6f64,
32'h68697073,
32'h68696e74,
32'h68657273,
32'h68657264,
32'h68657262,
32'h68656d70,
32'h6865656c,
32'h6865636b,
32'h68617473,
32'h68617468,
32'h68617368,
32'h68616c6f,
32'h6861636b,
32'h67757275,
32'h67756c66,
32'h676f776e,
32'h676f6174,
32'h676c6f77,
32'h67656d73,
32'h67617a65,
32'h67617073,
32'h66757365,
32'h66757279,
32'h66726f67,
32'h666f7274,
32'h666f726b,
32'h666f6f6c,
32'h666f6e64,
32'h666f6c6b,
32'h666f6c64,
32'h666f696c,
32'h666c6970,
32'h666c6578,
32'h666c6577,
32'h666c6564,
32'h66697374,
32'h66656174,
32'h66617473,
32'h66617265,
32'h66616465,
32'h6575726f,
32'h6563686f,
32'h65617473,
32'h6561726c,
32'h64756d70,
32'h64756d62,
32'h64756c6c,
32'h64756465,
32'h64756374,
32'h6475636b,
32'h646f7473,
32'h646f6f6d,
32'h646f6d65,
32'h646f6c6c,
32'h646f6373,
32'h646f636b,
32'h64697665,
32'h64696573,
32'h64696365,
32'h6469616c,
32'h64656564,
32'h64656166,
32'h6461776e,
32'h64617368,
32'h64617265,
32'h64616d70,
32'h64616d6e,
32'h63757265,
32'h63756c74,
32'h63756573,
32'h63756273,
32'h63756265,
32'h63726162,
32'h636f7a79,
32'h636f7773,
32'h636f7665,
32'h636f7073,
32'h636f7065,
32'h636f6e65,
32'h636f6b65,
32'h636f696c,
32'h636f636b,
32'h636c7565,
32'h636c616e,
32'h63686f70,
32'h6368696e,
32'h63686963,
32'h63686577,
32'h63617665,
32'h63617262,
32'h63616e73,
32'h63616e65,
32'h63616c6d,
32'h63616c66,
32'h63616765,
32'h63616665,
32'h62757973,
32'h62757474,
32'h62757368,
32'h62756d70,
32'h62756c6c,
32'h62756c62,
32'h62756473,
32'h6275636b,
32'h62726577,
32'h626f7574,
32'h626f7265,
32'h626f6f6d,
32'h626f696c,
32'h626c6577,
32'h626c6168,
32'h62697465,
32'h62696e64,
32'h62696473,
32'h62696173,
32'h62656e74,
32'h62656e64,
32'h62656c6c,
32'h62656573,
32'h6265616e,
32'h6265616d,
32'h62656164,
32'h62617473,
32'h6261726e,
32'h6261726b,
32'h62617265,
32'h62616e67,
32'h62616974,
32'h6261696c,
32'h61786c65,
32'h61766964,
32'h61757261,
32'h61756e74,
32'h61746f70,
32'h61746f6d,
32'h61726368,
32'h616e7473,
32'h616e7469,
32'h616d7073,
32'h616d6d6f,
32'h616d6964,
32'h616d656e,
32'h616c6c79,
32'h616c6173,
32'h616b696e,
32'h61676564,
32'h61637265,
32'h61636e65,
32'h7a65726f,
32'h796f6761,
32'h77726170,
32'h776f726e,
32'h776f7265,
32'h77697365,
32'h77696e73,
32'h77696e67,
32'h77617368,
32'h77616b65,
32'h77616765,
32'h76696365,
32'h756e746f,
32'h75676c79,
32'h7477696e,
32'h74756e65,
32'h746f7973,
32'h74697265,
32'h74696c6c,
32'h74696c65,
32'h74696572,
32'h74696564,
32'h74686f75,
32'h74656e74,
32'h7465656e,
32'h74616c65,
32'h7461696c,
32'h74616773,
32'h73796e63,
32'h73756974,
32'h73746972,
32'h7374656d,
32'h7370616d,
32'h736f7570,
32'h736f6e73,
32'h736f6c6f,
32'h736f6c65,
32'h736f6461,
32'h736f6170,
32'h736c6f74,
32'h736b6970,
32'h73697473,
32'h73696e67,
32'h73686f65,
32'h73686974,
32'h7365616c,
32'h7363616e,
32'h73616b65,
32'h726f7773,
32'h726f7365,
32'h726f7065,
32'h72656e74,
32'h72616e6b,
32'h7261696c,
32'h7261636b,
32'h71756974,
32'h70726f73,
32'h70726570,
32'h70726179,
32'h706f7572,
32'h706f6c6c,
32'h706f6c65,
32'h706c7567,
32'h706c6f74,
32'h70697065,
32'h70696e73,
32'h70657473,
32'h70617973,
32'h70616c6d,
32'h70616473,
32'h6f776e73,
32'h6f72616c,
32'h6f6b6179,
32'h6f696c73,
32'h6f646473,
32'h6e757473,
32'h6e6f6465,
32'h6e656174,
32'h6e617679,
32'h6e61696c,
32'h6d6f6f64,
32'h6d696e69,
32'h6d696c6c,
32'h6d696c64,
32'h6d657373,
32'h6d657368,
32'h6d657265,
32'h6d61736b,
32'h6d616c6c,
32'h6c6f636b,
32'h6c697073,
32'h6c696674,
32'h6c696573,
32'h6c656166,
32'h6c61776e,
32'h6b6e6565,
32'h6b697473,
32'h6b69636b,
32'h6b65656e,
32'h6a757279,
32'h6a6f6b65,
32'h6a617a7a,
32'h6a61696c,
32'h686f7365,
32'h686f6f6b,
32'h68697473,
32'h68697265,
32'h68696b65,
32'h68696465,
32'h6865616c,
32'h6861726d,
32'h67756e73,
32'h67726970,
32'h67726964,
32'h67726579,
32'h67726179,
32'h676c7565,
32'h67656e65,
32'h67617465,
32'h67616e67,
32'h666f6e74,
32'h666f616d,
32'h66617465,
32'h66616d65,
32'h66616b65,
32'h65786974,
32'h6576696c,
32'h65706963,
32'h65617273,
32'h64756b65,
32'h6472756d,
32'h64726577,
32'h64726167,
32'h6469736b,
32'h64697363,
32'h64697274,
32'h64656e79,
32'h64656d6f,
32'h64656572,
32'h64656172,
32'h63757473,
32'h63757073,
32'h63726f70,
32'h63726170,
32'h636f726e,
32'h636f7264,
32'h636f6e73,
32'h636f696e,
32'h636f6174,
32'h636f616c,
32'h636c6970,
32'h636c6179,
32'h63686970,
32'h63686566,
32'h63686174,
32'h63617274,
32'h63617073,
32'h6275726e,
32'h62756c6b,
32'h62756773,
32'h626f6f74,
32'h626f6e64,
32'h626f6d62,
32'h626f6c74,
32'h626f6c64,
32'h626c6f77,
32'h62697473,
32'h62657461,
32'h62656566,
32'h62656473,
32'h62656172,
32'h62617468,
32'h62617373,
32'h62616b65,
32'h61786973,
32'h61736b73,
32'h61696d73,
32'h61696473,
32'h7a6f6e65,
32'h796f7572,
32'h79656172,
32'h79656168,
32'h79617264,
32'h776f726b,
32'h776f7264,
32'h776f6f64,
32'h77697468,
32'h77697368,
32'h77697265,
32'h77696e65,
32'h77696e64,
32'h77696c6c,
32'h77696c64,
32'h77696665,
32'h77696465,
32'h77686f6d,
32'h7768656e,
32'h77686174,
32'h77657374,
32'h77657265,
32'h77656e74,
32'h77656c6c,
32'h7765656b,
32'h77656172,
32'h7765616b,
32'h77617973,
32'h77617665,
32'h77617273,
32'h7761726d,
32'h77616e74,
32'h77616c6c,
32'h77616c6b,
32'h77616974,
32'h766f7465,
32'h76697361,
32'h76696577,
32'h76657279,
32'h76617374,
32'h76617279,
32'h75736573,
32'h75736572,
32'h75736564,
32'h75706f6e,
32'h756e6974,
32'h74797065,
32'h7475726e,
32'h74756265,
32'h74726970,
32'h74726565,
32'h746f776e,
32'h746f7572,
32'h746f6f6c,
32'h746f6f6b,
32'h746f6e65,
32'h746f6c64,
32'h74697073,
32'h74696e79,
32'h74696d65,
32'h74687573,
32'h74686973,
32'h7468696e,
32'h74686579,
32'h7468656e,
32'h7468656d,
32'h74686174,
32'h7468616e,
32'h74657874,
32'h74657374,
32'h7465726d,
32'h74656e64,
32'h74656c6c,
32'h74656368,
32'h7465616d,
32'h7461736b,
32'h74617065,
32'h74616e6b,
32'h74616c6c,
32'h74616c6b,
32'h74616b65,
32'h73757265,
32'h73756368,
32'h73746f70,
32'h73746570,
32'h73746179,
32'h73746172,
32'h73706f74,
32'h736f756c,
32'h736f7274,
32'h736f6f6e,
32'h736f6e67,
32'h736f6d65,
32'h736f6c64,
32'h736f696c,
32'h736f6674,
32'h736e6f77,
32'h736c6f77,
32'h736b696e,
32'h73697a65,
32'h73697465,
32'h7369676e,
32'h73696465,
32'h7369636b,
32'h73687574,
32'h73686f77,
32'h73686f74,
32'h73686f70,
32'h73686970,
32'h73657473,
32'h73656e74,
32'h73656e64,
32'h73656c6c,
32'h73656c66,
32'h73656573,
32'h7365656e,
32'h7365656d,
32'h7365656b,
32'h73656564,
32'h73656174,
32'h73617973,
32'h73617665,
32'h73616e64,
32'h73616d65,
32'h73616c74,
32'h73616c65,
32'h73616964,
32'h73616665,
32'h72756e73,
32'h72756c65,
32'h726f6f74,
32'h726f6f6d,
32'h726f6f66,
32'h726f6c6c,
32'h726f6c65,
32'h726f636b,
32'h726f6164,
32'h7269736b,
32'h72697365,
32'h72696e67,
32'h72696465,
32'h72696368,
32'h72696365,
32'h72657374,
32'h72656c79,
32'h72656172,
32'h7265616c,
32'h72656164,
32'h72617465,
32'h72617265,
32'h7261696e,
32'h72616365,
32'h70757473,
32'h70757368,
32'h70757265,
32'h70756d70,
32'h70756c6c,
32'h706f7374,
32'h706f7274,
32'h706f6f72,
32'h706f6f6c,
32'h706c7573,
32'h706c6179,
32'h706c616e,
32'h70696e6b,
32'h7069636b,
32'h7065616b,
32'h70617468,
32'h70617374,
32'h70617373,
32'h70617274,
32'h7061726b,
32'h70616972,
32'h7061696e,
32'h70616964,
32'h70616765,
32'h7061636b,
32'h70616365,
32'h6f766572,
32'h6f76656e,
32'h6f70656e,
32'h6f6e746f,
32'h6f6e6c79,
32'h6f6e6573,
32'h6f6e6365,
32'h6e6f7465,
32'h6e6f7365,
32'h6e6f6e65,
32'h6e696e65,
32'h6e696365,
32'h6e657874,
32'h6e657773,
32'h6e656564,
32'h6e65636b,
32'h6e656172,
32'h6e616d65,
32'h6d757374,
32'h6d756368,
32'h6d6f7665,
32'h6d6f7374,
32'h6d6f7265,
32'h6d6f6f6e,
32'h6d6f6465,
32'h6d697373,
32'h6d696e65,
32'h6d696e64,
32'h6d696c6b,
32'h6d696c65,
32'h6d656e75,
32'h6d656574,
32'h6d656174,
32'h6d65616e,
32'h6d65616c,
32'h6d617468,
32'h6d617373,
32'h6d61726b,
32'h6d617073,
32'h6d616e79,
32'h6d616c65,
32'h6d616b65,
32'h6d61696e,
32'h6d61696c,
32'h6d616465,
32'h6c75636b,
32'h6c6f7665,
32'h6c6f7473,
32'h6c6f7374,
32'h6c6f7373,
32'h6c6f7365,
32'h6c6f7264,
32'h6c6f6f70,
32'h6c6f6f6b,
32'h6c6f6e67,
32'h6c6f676f,
32'h6c6f616e,
32'h6c6f6164,
32'h6c697665,
32'h6c697374,
32'h6c696e6b,
32'h6c696e65,
32'h6c696b65,
32'h6c696665,
32'h6c657373,
32'h6c656e73,
32'h6c656773,
32'h6c656674,
32'h6c656164,
32'h6c617773,
32'h6c617465,
32'h6c617374,
32'h6c616e65,
32'h6c616e64,
32'h6c616b65,
32'h6c616964,
32'h6c616479,
32'h6c61636b,
32'h6b6e6f77,
32'h6b6e6577,
32'h6b696e67,
32'h6b696e64,
32'h6b696c6c,
32'h6b696473,
32'h6b657973,
32'h6b657074,
32'h6b656570,
32'h6a757374,
32'h6a756d70,
32'h6a6f696e,
32'h6a6f6273,
32'h6974656d,
32'h69726f6e,
32'h696e746f,
32'h696e666f,
32'h696e6368,
32'h69646561,
32'h69636f6e,
32'h68757274,
32'h68756765,
32'h686f7572,
32'h686f7374,
32'h686f7065,
32'h686f6d65,
32'h686f6c79,
32'h686f6c65,
32'h686f6c64,
32'h68696c6c,
32'h68696768,
32'h6865726f,
32'h68657265,
32'h68656c70,
32'h68656c6c,
32'h68656c64,
32'h68656174,
32'h68656172,
32'h68656164,
32'h68617665,
32'h68617465,
32'h68617264,
32'h68616e67,
32'h68616e64,
32'h68616c6c,
32'h68616c66,
32'h68616972,
32'h67757973,
32'h67726f77,
32'h67726577,
32'h67726162,
32'h676f6f64,
32'h676f6e65,
32'h676f6c66,
32'h676f6c64,
32'h676f6573,
32'h676f6473,
32'h676f616c,
32'h676c6164,
32'h67697665,
32'h6769726c,
32'h67696674,
32'h67657473,
32'h67656172,
32'h67617665,
32'h67616d65,
32'h6761696e,
32'h66756e64,
32'h66756c6c,
32'h6675656c,
32'h66726f6d,
32'h66726565,
32'h666f7572,
32'h666f726d,
32'h666f6f74,
32'h666f6f64,
32'h666c6f77,
32'h666c6174,
32'h666c6167,
32'h66697665,
32'h66697473,
32'h66697368,
32'h6669726d,
32'h66697265,
32'h66696e65,
32'h66696e64,
32'h66696c6d,
32'h66696c6c,
32'h66696c65,
32'h66656c74,
32'h66656c6c,
32'h66656574,
32'h66656573,
32'h6665656c,
32'h66656564,
32'h66656172,
32'h66617374,
32'h6661726d,
32'h66616e73,
32'h66616c6c,
32'h66616972,
32'h6661696c,
32'h66616374,
32'h66616365,
32'h65796573,
32'h6578616d,
32'h65766572,
32'h6576656e,
32'h656e6473,
32'h656c7365,
32'h65676773,
32'h65646974,
32'h65646765,
32'h65617379,
32'h65617374,
32'h65617365,
32'h6561726e,
32'h65616368,
32'h64757479,
32'h64757374,
32'h6475616c,
32'h64727567,
32'h64726f70,
32'h64726177,
32'h646f776e,
32'h646f7365,
32'h646f6f72,
32'h646f6e65,
32'h646f6773,
32'h646f6573,
32'h64697368,
32'h64696574,
32'h64696564,
32'h6465736b,
32'h64656570,
32'h6465636b,
32'h64656274,
32'h6465616c,
32'h64656164,
32'h64617973,
32'h64617465,
32'h64617461,
32'h6461726b,
32'h63757465,
32'h63726577,
32'h636f7374,
32'h636f7265,
32'h636f7079,
32'h636f6f6c,
32'h636f6f6b,
32'h636f6d65,
32'h636f6c64,
32'h636f6465,
32'h636c7562,
32'h63697479,
32'h63656e74,
32'h63656c6c,
32'h63617473,
32'h63617374,
32'h63617368,
32'h63617365,
32'h63617273,
32'h63617265,
32'h63617264,
32'h63616d70,
32'h63616d65,
32'h63616c6c,
32'h63616b65,
32'h62757379,
32'h626f7973,
32'h626f776c,
32'h626f7468,
32'h626f7373,
32'h626f726e,
32'h626f6f6b,
32'h626f6e65,
32'h626f6479,
32'h626f6174,
32'h626c7565,
32'h626c6f67,
32'h62697264,
32'h62696c6c,
32'h62696b65,
32'h62657374,
32'h62656c74,
32'h62656572,
32'h6265656e,
32'h62656174,
32'h62617365,
32'h62617273,
32'h62616e6b,
32'h62616e64,
32'h62616c6c,
32'h62616773,
32'h6261636b,
32'h62616279,
32'h61776179,
32'h6175746f,
32'h61727473,
32'h61726d79,
32'h61726d73,
32'h61726561,
32'h61707073,
32'h616c736f,
32'h61676573,
32'h61646473,
32'h61637473,
32'h61636964,
32'h61626c65
};

localparam bit [7:0] MAP_SHORT [0:31] = '{
    8'h65, 8'h20, 8'h6b, 8'h69, 8'h6e, 8'h67, 8'h6d, 8'h6f, 
    8'h6c, 8'h74, 8'h61, 8'h72, 8'h73, 8'h68, 8'h64, 8'h75, 
    8'h77, 8'h66, 8'h63, 8'h79, 8'h70, 8'h62, 8'h76, 8'h6a, 
    8'h78, 8'h71, 8'h7a, 8'h2c, 8'h2e, 8'h5f, 8'h3f, 8'h21
};

localparam bit [7:0] MAP_LONG [0:63] = '{
    8'h65, 8'h20, 8'h74, 8'h61, 8'h72, 8'h69, 8'h6f, 8'h6e, 
    8'h73, 8'h68, 8'h64, 8'h6c, 8'h75, 8'h77, 8'h6d, 8'h66, 
    8'h63, 8'h67, 8'h79, 8'h70, 8'h62, 8'h6b, 8'h76, 8'h6a, 
    8'h78, 8'h71, 8'h7a, 8'h2c, 8'h2e, 8'h3f, 8'h21, 8'h45, 
    8'h54, 8'h41, 8'h52, 8'h49, 8'h4f, 8'h4e, 8'h53, 8'h48, 
    8'h44, 8'h4c, 8'h55, 8'h57, 8'h4d, 8'h46, 8'h43, 8'h47, 
    8'h59, 8'h50, 8'h42, 8'h4b, 8'h4a, 8'h58, 8'h30, 8'h31, 
    8'h32, 8'h33, 8'h34, 8'h35, 8'h36, 8'h37, 8'h38, 8'h39
};

reg [11:0] counter_dict_reg, counter_dict_next;
reg [29:0] counter_short_reg, counter_short_next;
reg [35:0] counter_long_reg, counter_long_next;

localparam STATE_SIZE = 2;
localparam [STATE_SIZE-1:0] dict = 2'h0,
                            short = 2'h1,
                            long = 2'h2,
                            fini = 2'h3;


reg [STATE_SIZE-1:0] state_reg, state_next;

reg [47:0] key_reg, key_next;

reg [33:0] start_reg, start_next;
reg [33:0] valid_reg, valid_next;
reg rdy_reg, rdy_next;

reg [5:0] decryptor_counter_reg, decryptor_counter_next;

reg [47:0] final_key_reg, final_key_next;

assign valid = valid_reg > 0;
assign rdy = rdy_reg;
assign key_out = final_key_reg;

wire [0:33] [47:0] temp_key;

always@(posedge clk, posedge rst) begin
    if(rst) begin
        counter_dict_reg <= 0;
        counter_short_reg <= 0;
        counter_long_reg <= 0;
        
        decryptor_counter_reg <= 0;
        valid_reg <= 0;
        start_reg <= 0;
        rdy_reg <= 0;
        
        final_key_reg <= 0;
        
        key_reg <= 0;
        state_reg <= dict;
    end else begin
        counter_dict_reg <= counter_dict_next;
        counter_short_reg <= counter_short_next;
        counter_long_reg <= counter_long_next; 
        
        decryptor_counter_reg <= decryptor_counter_next;
        valid_reg <= valid_next;
        start_reg <= start_next;
        rdy_reg <= rdy_next;
        
        final_key_reg <= final_key_next;
        
        key_reg <= key_next;
        state_reg <= state_next;
    end
end

always@(*) begin
    case(state_reg) 
        dict: state_next = valid ? fini : counter_dict_next > DICT4_SIZE ? short : dict;
        short: state_next = valid ? fini : counter_short_next == 0 ? long : short;
        long: state_next = valid || counter_long_next == 0 ? fini : long;
        fini: state_next = fini;
    endcase
end

always@(*) begin
    counter_dict_next = 0;
    counter_short_next = 0;
    counter_long_next = 0;
    key_next = 0;
    rdy_next = 0;
    final_key_next = final_key_reg;
    
    if(decryptor_counter_reg >= 34) 
        decryptor_counter_next = 0;
    else 
        decryptor_counter_next = decryptor_counter_reg + 1'b1;
        
    start_next = 1 << decryptor_counter_reg;
    
    case(state_reg) 
        dict: begin
            counter_dict_next = counter_dict_reg + 1'b1;
            key_next = {"e ", DICT4[counter_dict_reg]};
        end
        short: begin
            counter_short_next = counter_short_reg + 1'b1;
            key_next = {
                MAP_SHORT[counter_short_reg[29:25]],
                MAP_SHORT[counter_short_reg[24:20]],
                MAP_SHORT[counter_short_reg[19:15]],
                MAP_SHORT[counter_short_reg[14:10]],
                MAP_SHORT[counter_short_reg[9:5]],
                MAP_SHORT[counter_short_reg[4:0]]
            };
        end
        long: begin
            counter_long_next = counter_long_reg + 1'b1;
            key_next = {
                MAP_LONG[counter_long_reg[35:30]],
                MAP_LONG[counter_long_reg[29:24]],
                MAP_LONG[counter_long_reg[23:18]],
                MAP_LONG[counter_long_reg[17:12]],
                MAP_LONG[counter_long_reg[11:6]],
                MAP_LONG[counter_long_reg[5:0]]
            };
        end
        fini: begin
            rdy_next = 1;
            if(!rdy_reg)
                final_key_next = temp_key[33];
        end
    endcase
end

genvar i;

generate
    wire [47:0] key_out_gen;
    
    for (i = 0; i < 34; i = i + 1) begin : generate_block_identifier
        wire [47:0] key_out_tmp;
         
        tea_asmd d0 (
            .clk(clk),
            .rst(rst),
            .ena(ena),
            .start(start_reg[i]),
            .data(data),
            .key(key_next),
            .key_out(key_out_tmp),
            .valid(valid_next[i])
        );
        
        if(i > 0) begin
            assign temp_key[i] = temp_key[i - 1] | ({48{valid_reg[i]}} & key_out_tmp);
        end else begin
            assign temp_key[i] = ({48{valid_reg[i]}} & key_out_tmp);
        end
    end
endgenerate

endmodule
